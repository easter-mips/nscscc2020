`ifndef DCACHE_DEFS_SVH
`define DCACHE_DEFS_SVH

typedef logic[31:0] Data;
typedef logic[31:0] Addr;

typedef Data[7:0] WayBankData;

`endif